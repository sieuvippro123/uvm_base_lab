interface vip_clkrst_intf;
    //-------------------------------------------------------------------------
    //  Signals
    //-------------------------------------------------------------------------
    logic   clk     ;   //  Clock
    logic   resetn  ;   //  Asynchronous active low reset

    //-------------------------------------------------------------------------
    //  Modport
    //-------------------------------------------------------------------------
    modport TEST(
        output  clk     ,
        output  resetn
    );

endinterface
