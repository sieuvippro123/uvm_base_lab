interface vip_sig_mnt_intf();
    //-------------------------------------------------------------------------
    //  Interface Signals
    //-------------------------------------------------------------------------
    logic       mnt_sig ;

    //-------------------------------------------------------------------------
    //  Modport
    //-------------------------------------------------------------------------
    modport TEST(
        input   mnt_sig
    );

endinterface
